set_property PACKAGE_PIN V2 [get_ports {num2[0]}]
set_property IOSTANDARD LVCMOS33 [get_ports {num2[0]}]
set_property PACKAGE_PIN T3 [get_ports {num2[1]}]
set_property IOSTANDARD LVCMOS33 [get_ports {num2[1]}]
set_property PACKAGE_PIN T2 [get_ports {num2[2]}]
set_property IOSTANDARD LVCMOS33 [get_ports {num2[2]}]
set_property PACKAGE_PIN R3 [get_ports {num2[3]}]
set_property IOSTANDARD LVCMOS33 [get_ports {num2[3]}]
set_property PACKAGE_PIN W2 [get_ports {num1[0]}]
set_property IOSTANDARD LVCMOS33 [get_ports {num1[0]}]
set_property PACKAGE_PIN U1 [get_ports {num1[1]}]
set_property IOSTANDARD LVCMOS33 [get_ports {num1[1]}]
set_property PACKAGE_PIN T1 [get_ports {num1[2]}]
set_property IOSTANDARD LVCMOS33 [get_ports {num1[2]}]
set_property PACKAGE_PIN R2 [get_ports {num1[3]}]
set_property IOSTANDARD LVCMOS33 [get_ports {num1[3]}]

set_property PACKAGE_PIN V17 [get_ports {sel[0]}]
set_property IOSTANDARD LVCMOS33 [get_ports {sel[0]}]
set_property PACKAGE_PIN V16 [get_ports {sel[1]}]
set_property IOSTANDARD LVCMOS33 [get_ports {sel[1]}]
set_property PACKAGE_PIN W16 [get_ports {sel[2]}]
set_property IOSTANDARD LVCMOS33 [get_ports {sel[2]}]

set_property PACKAGE_PIN P3 [get_ports {func_o[0]}]
set_property IOSTANDARD LVCMOS33 [get_ports {func_o[0]}]
set_property PACKAGE_PIN N3 [get_ports {func_o[1]}]
set_property IOSTANDARD LVCMOS33 [get_ports {func_o[1]}]
set_property PACKAGE_PIN P1 [get_ports {func_o[2]}]
set_property IOSTANDARD LVCMOS33 [get_ports {func_o[2]}]
set_property PACKAGE_PIN L1 [get_ports {func_o[3]}]
set_property IOSTANDARD LVCMOS33 [get_ports {func_o[3]}]

set_property PACKAGE_PIN U16 [get_ports {overflow}]
set_property IOSTANDARD LVCMOS33 [get_ports {overflow}]
